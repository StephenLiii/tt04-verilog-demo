`default_nettype none
`timescale 1ns / 1ps

module rom_sprite_cat (
    input wire [9:0] addr,
    output reg [3:0] data
);

always @(*) begin
    case (addr)
        10'd0: data = 4'h6;
        10'd1: data = 4'h6;
        10'd2: data = 4'h6;
        10'd3: data = 4'h6;
        10'd4: data = 4'h6;
        10'd5: data = 4'h6;
        10'd6: data = 4'h6;
        10'd7: data = 4'h6;
        10'd8: data = 4'h6;
        10'd9: data = 4'h6;
        10'd10: data = 4'h6;
        10'd11: data = 4'h6;
        10'd12: data = 4'h6;
        10'd13: data = 4'h6;
        10'd14: data = 4'h6;
        10'd15: data = 4'h6;
        10'd16: data = 4'h6;
        10'd17: data = 4'h6;
        10'd18: data = 4'h6;
        10'd19: data = 4'h6;
        10'd20: data = 4'h6;
        10'd21: data = 4'h6;
        10'd22: data = 4'h6;
        10'd23: data = 4'h6;
        10'd24: data = 4'h6;
        10'd25: data = 4'h6;
        10'd26: data = 4'h6;
        10'd27: data = 4'h6;
        10'd28: data = 4'h6;
        10'd29: data = 4'h6;
        10'd30: data = 4'h6;
        10'd31: data = 4'h6;
        10'd32: data = 4'h6;
        10'd33: data = 4'h6;
        10'd34: data = 4'h6;
        10'd35: data = 4'h6;
        10'd36: data = 4'h6;
        10'd37: data = 4'h6;
        10'd38: data = 4'h6;
        10'd39: data = 4'h6;
        10'd40: data = 4'h6;
        10'd41: data = 4'h6;
        10'd42: data = 4'h6;
        10'd43: data = 4'h6;
        10'd44: data = 4'h6;
        10'd45: data = 4'h6;
        10'd46: data = 4'h6;
        10'd47: data = 4'h6;
        10'd48: data = 4'h6;
        10'd49: data = 4'h6;
        10'd50: data = 4'h6;
        10'd51: data = 4'h6;
        10'd52: data = 4'h6;
        10'd53: data = 4'h6;
        10'd54: data = 4'h6;
        10'd55: data = 4'h6;
        10'd56: data = 4'h6;
        10'd57: data = 4'h6;
        10'd58: data = 4'h6;
        10'd59: data = 4'h6;
        10'd60: data = 4'h6;
        10'd61: data = 4'h6;
        10'd62: data = 4'h6;
        10'd63: data = 4'h6;
        10'd64: data = 4'h6;
        10'd65: data = 4'h6;
        10'd66: data = 4'h6;
        10'd67: data = 4'h6;
        10'd68: data = 4'h6;
        10'd69: data = 4'h6;
        10'd70: data = 4'h6;
        10'd71: data = 4'h6;
        10'd72: data = 4'h6;
        10'd73: data = 4'h6;
        10'd74: data = 4'h6;
        10'd75: data = 4'h6;
        10'd76: data = 4'h6;
        10'd77: data = 4'h6;
        10'd78: data = 4'h6;
        10'd79: data = 4'h6;
        10'd80: data = 4'h6;
        10'd81: data = 4'h6;
        10'd82: data = 4'h6;
        10'd83: data = 4'h6;
        10'd84: data = 4'h6;
        10'd85: data = 4'h6;
        10'd86: data = 4'h6;
        10'd87: data = 4'h6;
        10'd88: data = 4'h6;
        10'd89: data = 4'h6;
        10'd90: data = 4'h6;
        10'd91: data = 4'h6;
        10'd92: data = 4'h6;
        10'd93: data = 4'h6;
        10'd94: data = 4'h6;
        10'd95: data = 4'h5;
        10'd96: data = 4'h6;
        10'd97: data = 4'h6;
        10'd98: data = 4'h6;
        10'd99: data = 4'h6;
                10'd100: data = 4'h6;
        10'd101: data = 4'h6;
        10'd102: data = 4'h6;
        10'd103: data = 4'h6;
        10'd104: data = 4'h6;
        10'd105: data = 4'h6;
        10'd106: data = 4'h6;
        10'd107: data = 4'h6;
        10'd108: data = 4'h6;
        10'd109: data = 4'h6;
        10'd110: data = 4'h6;
        10'd111: data = 4'h6;
        10'd112: data = 4'h6;
        10'd113: data = 4'h6;
        10'd114: data = 4'h6;
        10'd115: data = 4'h6;
        10'd116: data = 4'h6;
        10'd117: data = 4'h6;
        10'd118: data = 4'h6;
        10'd119: data = 4'h6;
        10'd120: data = 4'h6;
        10'd121: data = 4'h6;
        10'd122: data = 4'h6;
        10'd123: data = 4'h6;
        10'd124: data = 4'h6;
        10'd125: data = 4'h5;
        10'd126: data = 4'h6;
        10'd127: data = 4'h6;
        10'd128: data = 4'h6;
        10'd129: data = 4'h6;
        10'd130: data = 4'h5;
        10'd131: data = 4'h1;
        10'd132: data = 4'h5;
        10'd133: data = 4'h6;
        10'd134: data = 4'h6;
        10'd135: data = 4'h6;
        10'd136: data = 4'h6;
        10'd137: data = 4'h6;
        10'd138: data = 4'h6;
        10'd139: data = 4'h5;
        10'd140: data = 4'h1;
        10'd141: data = 4'h5;
        10'd142: data = 4'h6;
        10'd143: data = 4'h6;
        10'd144: data = 4'h6;
        10'd145: data = 4'h6;
        10'd146: data = 4'h5;
        10'd147: data = 4'h1;
        10'd148: data = 4'h5;
        10'd149: data = 4'h6;
        10'd150: data = 4'h6;
        10'd151: data = 4'h6;
        10'd152: data = 4'h6;
        10'd153: data = 4'h6;
        10'd154: data = 4'h6;
        10'd155: data = 4'h5;
        10'd156: data = 4'h1;
        10'd157: data = 4'h1;
        10'd158: data = 4'h5;
        10'd159: data = 4'h5;
        10'd160: data = 4'h5;
        10'd161: data = 4'h5;
        10'd162: data = 4'h5;
        10'd163: data = 4'h5;
        10'd164: data = 4'h1;
        10'd165: data = 4'h0;
        10'd166: data = 4'h5;
        10'd167: data = 4'h6;
        10'd168: data = 4'h6;
        10'd169: data = 4'h6;
        10'd170: data = 4'h6;
        10'd171: data = 4'h5;
        10'd172: data = 4'h1;
        10'd173: data = 4'h0;
        10'd174: data = 4'h5;
        10'd175: data = 4'h6;
        10'd176: data = 4'h6;
        10'd177: data = 4'h6;
        10'd178: data = 4'h6;
        10'd179: data = 4'h6;
        10'd180: data = 4'h6;
        10'd181: data = 4'h5;
        10'd182: data = 4'h1;
        10'd183: data = 4'h1;
        10'd184: data = 4'h1;
        10'd185: data = 4'h1;
        10'd186: data = 4'h1;
        10'd187: data = 4'h1;
        10'd188: data = 4'h1;
        10'd189: data = 4'h1;
        10'd190: data = 4'h1;
        10'd191: data = 4'h1;
        10'd192: data = 4'h5;
        10'd193: data = 4'h6;
        10'd194: data = 4'h6;
        10'd195: data = 4'h6;
        10'd196: data = 4'h5;
        10'd197: data = 4'h1;
        10'd198: data = 4'h0;
        10'd199: data = 4'h5;
                10'd200: data = 4'h6;
        10'd201: data = 4'h6;
        10'd202: data = 4'h6;
        10'd203: data = 4'h6;
        10'd204: data = 4'h5;
        10'd205: data = 4'h1;
        10'd206: data = 4'h0;
        10'd207: data = 4'h5;
        10'd208: data = 4'h6;
        10'd209: data = 4'h6;
        10'd210: data = 4'h6;
        10'd211: data = 4'h6;
        10'd212: data = 4'h5;
        10'd213: data = 4'h1;
        10'd214: data = 4'h1;
        10'd215: data = 4'h5;
        10'd216: data = 4'h5;
        10'd217: data = 4'h5;
        10'd218: data = 4'h5;
        10'd219: data = 4'h5;
        10'd220: data = 4'h5;
        10'd221: data = 4'h1;
        10'd222: data = 4'h0;
        10'd223: data = 4'h5;
        10'd224: data = 4'h6;
        10'd225: data = 4'h5;
        10'd226: data = 4'h1;
        10'd227: data = 4'h0;
        10'd228: data = 4'h5;
        10'd229: data = 4'h6;
        10'd230: data = 4'h5;
        10'd231: data = 4'h1;
        10'd232: data = 4'h0;
        10'd233: data = 4'h5;
        10'd234: data = 4'h5;
        10'd235: data = 4'h5;
        10'd236: data = 4'h5;
        10'd237: data = 4'h5;
        10'd238: data = 4'h0;
        10'd239: data = 4'h5;
        10'd240: data = 4'h5;
        10'd241: data = 4'h5;
        10'd242: data = 4'h5;
        10'd243: data = 4'h0;
        10'd244: data = 4'h5;
        10'd245: data = 4'h5;
        10'd246: data = 4'h5;
        10'd247: data = 4'h5;
        10'd248: data = 4'h5;
        10'd249: data = 4'h5;
        10'd250: data = 4'h5;
        10'd251: data = 4'h5;
        10'd252: data = 4'h5;
        10'd253: data = 4'h5;
        10'd254: data = 4'h5;
        10'd255: data = 4'h5;
        10'd256: data = 4'h5;
        10'd257: data = 4'h5;
        10'd258: data = 4'h5;
        10'd259: data = 4'h5;
        10'd260: data = 4'h5;
        10'd261: data = 4'h5;
        10'd262: data = 4'h5;
        10'd263: data = 4'h5;
        10'd264: data = 4'h5;
        10'd265: data = 4'h5;
        10'd266: data = 4'h5;
        10'd267: data = 4'h5;
        10'd268: data = 4'h5;
        10'd269: data = 4'h5;
        10'd270: data = 4'h5;
        10'd271: data = 4'h5;
        10'd272: data = 4'h5;
        10'd273: data = 4'h5;
        10'd274: data = 4'h5;
        10'd275: data = 4'h5;
        10'd276: data = 4'h5;
        10'd277: data = 4'h5;
        10'd278: data = 4'h5;
        10'd279: data = 4'h5;
        10'd280: data = 4'h5;
        10'd281: data = 4'h5;
        10'd282: data = 4'h5;
        10'd283: data = 4'h5;
        10'd284: data = 4'h5;
        10'd285: data = 4'h5;
        10'd286: data = 4'h5;
        10'd287: data = 4'h5;
        10'd288: data = 4'h5;
        10'd289: data = 4'h5;
        10'd290: data = 4'h5;
        10'd291: data = 4'h5;
        10'd292: data = 4'h5;
        10'd293: data = 4'h5;
        10'd294: data = 4'h5;
        10'd295: data = 4'h5;
        10'd296: data = 4'h5;
        10'd297: data = 4'h5;
        10'd298: data = 4'h5;
        10'd299: data = 4'h5;
                10'd300: data = 4'h5;
        10'd301: data = 4'h1;
        10'd302: data = 4'h1;
        10'd303: data = 4'h5;
        10'd304: data = 4'h5;
        10'd305: data = 4'h1;
        10'd306: data = 4'h1;
        10'd307: data = 4'h5;
        10'd308: data = 4'h5;
        10'd309: data = 4'h1;
        10'd310: data = 4'h1;
        10'd311: data = 4'h5;
        10'd312: data = 4'h5;
        10'd313: data = 4'h1;
        10'd314: data = 4'h1;
        10'd315: data = 4'h5;
        10'd316: data = 4'h5;
        10'd317: data = 4'h5;
        10'd318: data = 4'h5;
        10'd319: data = 4'h5;
        10'd320: data = 4'h5;
        10'd321: data = 4'h1;
        10'd322: data = 4'h1;
        10'd323: data = 4'h5;
        10'd324: data = 4'h5;
        10'd325: data = 4'h5;
        10'd326: data = 4'h5;
        10'd327: data = 4'h5;
        10'd328: data = 4'h5;
        10'd329: data = 4'h1;
        10'd330: data = 4'h1;
        10'd331: data = 4'h5;
        10'd332: data = 4'h5;
        10'd333: data = 4'h5;
        10'd334: data = 4'h5;
        10'd335: data = 4'h5;
        10'd336: data = 4'h5;
        10'd337: data = 4'h5;
        10'd338: data = 4'h5;
        10'd339: data = 4'h5;
        10'd340: data = 4'h5;
        10'd341: data = 4'h5;
        10'd342: data = 4'h5;
        10'd343: data = 4'h5;
        10'd344: data = 4'h5;
        10'd345: data = 4'h5;
        10'd346: data = 4'h5;
        10'd347: data = 4'h5;
        10'd348: data = 4'h5;
        10'd349: data = 4'h5;
        10'd350: data = 4'h5;
        10'd351: data = 4'h5;
        10'd352: data = 4'h5;
        10'd353: data = 4'h5;
        10'd354: data = 4'h5;
        10'd355: data = 4'h5;
        10'd356: data = 4'h5;
        10'd357: data = 4'h5;
        10'd358: data = 4'h5;
        10'd359: data = 4'h5;
        10'd360: data = 4'h5;
        10'd361: data = 4'h5;
        10'd362: data = 4'h5;
        10'd363: data = 4'h5;
        10'd364: data = 4'h5;
        10'd365: data = 4'h5;
        10'd366: data = 4'h5;
        10'd367: data = 4'h5;
        10'd368: data = 4'h5;
        10'd369: data = 4'h5;
        10'd370: data = 4'h5;
        10'd371: data = 4'h5;
        10'd372: data = 4'h5;
        10'd373: data = 4'h5;
        10'd374: data = 4'h5;
        10'd375: data = 4'h5;
        10'd376: data = 4'h5;
        10'd377: data = 4'h5;
        10'd378: data = 4'h5;
        10'd379: data = 4'h5;
        10'd380: data = 4'h5;
        10'd381: data = 4'h5;
        10'd382: data = 4'h5;
        10'd383: data = 4'h5;
        10'd384: data = 4'h5;
        10'd385: data = 4'h5;
        10'd386: data = 4'h5;
        10'd387: data = 4'h5;
        10'd388: data = 4'h5;
        10'd389: data = 4'h5;
        10'd390: data = 4'h5;
        10'd391: data = 4'h5;
        10'd392: data = 4'h5;
        10'd393: data = 4'h5;
        10'd394: data = 4'h5;
        10'd395: data = 4'h5;
        10'd396: data = 4'h5;
        10'd397: data = 4'h5;
        10'd398: data = 4'h5;
        10'd399: data = 4'h5;
                10'd400: data = 4'h5;
        10'd401: data = 4'h5;
        10'd402: data = 4'h1;
        10'd403: data = 4'h1;
        10'd404: data = 4'h5;
        10'd405: data = 4'h5;
        10'd406: data = 4'h1;
        10'd407: data = 4'h1;
        10'd408: data = 4'h5;
        10'd409: data = 4'h5;
        10'd410: data = 4'h4;
        10'd411: data = 4'h4;
        10'd412: data = 4'h2;
        10'd413: data = 4'h1;
        10'd414: data = 4'h1;
        10'd415: data = 4'h1;
        10'd416: data = 4'h0;
        10'd417: data = 4'h5;
        10'd418: data = 4'h5;
        10'd419: data = 4'h5;
        10'd420: data = 4'h0;
        10'd421: data = 4'h5;
        10'd422: data = 4'h6;
        10'd423: data = 4'h6;
        10'd424: data = 4'h6;
        10'd425: data = 4'h6;
        10'd426: data = 4'h5;
        10'd427: data = 4'h5;
        10'd428: data = 4'h2;
        10'd429: data = 4'h2;
        10'd430: data = 4'h2;
        10'd431: data = 4'h2;
        10'd432: data = 4'h1;
        10'd433: data = 4'h0;
        10'd434: data = 4'h0;
        10'd435: data = 4'h1;
        10'd436: data = 4'h1;
        10'd437: data = 4'h3;
        10'd438: data = 4'h1;
        10'd439: data = 4'h0;
        10'd440: data = 4'h5;
        10'd441: data = 4'h6;
        10'd442: data = 4'h6;
        10'd443: data = 4'h6;
        10'd444: data = 4'h6;
        10'd445: data = 4'h6;
        10'd446: data = 4'h6;
        10'd447: data = 4'h5;
        10'd448: data = 4'h0;
        10'd449: data = 4'h0;
        10'd450: data = 4'h0;
        10'd451: data = 4'h0;
        10'd452: data = 4'h0;
        10'd453: data = 4'h0;
        10'd454: data = 4'h3;
        10'd455: data = 4'h1;
        10'd456: data = 4'h1;
        10'd457: data = 4'h3;
        10'd458: data = 4'h0;
        10'd459: data = 4'h5;
        10'd460: data = 4'h6;
        10'd461: data = 4'h6;
        10'd462: data = 4'h6;
        10'd463: data = 4'h6;
        10'd464: data = 4'h6;
        10'd465: data = 4'h6;
        10'd466: data = 4'h5;
        10'd467: data = 4'h1;
        10'd468: data = 4'h3;
        10'd469: data = 4'h1;
        10'd470: data = 4'h3;
        10'd471: data = 4'h1;
        10'd472: data = 4'h1;
        10'd473: data = 4'h3;
        10'd474: data = 4'h1;
        10'd475: data = 4'h1;
        10'd476: data = 4'h1;
        10'd477: data = 4'h0;
        10'd478: data = 4'h5;
        10'd479: data = 4'h6;
        10'd480: data = 4'h6;
        10'd481: data = 4'h6;
        10'd482: data = 4'h6;
        10'd483: data = 4'h6;
        10'd484: data = 4'h6;
        10'd485: data = 4'h5;
        10'd486: data = 4'h1;
        10'd487: data = 4'h3;
        10'd488: data = 4'h1;
        10'd489: data = 4'h3;
        10'd490: data = 4'h1;
        10'd491: data = 4'h1;
        10'd492: data = 4'h1;
        10'd493: data = 4'h1;
        10'd494: data = 4'h1;
        10'd495: data = 4'h5;
        10'd496: data = 4'h6;
        10'd497: data = 4'h6;
        10'd498: data = 4'h6;
        10'd499: data = 4'h6;
                10'd500: data = 4'h6;
        10'd501: data = 4'h6;
        10'd502: data = 4'h6;
        10'd503: data = 4'h5;
        10'd504: data = 4'h1;
        10'd505: data = 4'h1;
        10'd506: data = 4'h1;
        10'd507: data = 4'h1;
        10'd508: data = 4'h5;
        10'd509: data = 4'h5;
        10'd510: data = 4'h5;
        10'd511: data = 4'h1;
        10'd512: data = 4'h1;
        10'd513: data = 4'h1;
        10'd514: data = 4'h5;
        10'd515: data = 4'h6;
        10'd516: data = 4'h5;
        10'd517: data = 4'h1;
        10'd518: data = 4'h1;
        10'd519: data = 4'h1;
        10'd520: data = 4'h5;
        10'd521: data = 4'h6;
        10'd522: data = 4'h5;
        10'd523: data = 4'h1;
        10'd524: data = 4'h1;
        10'd525: data = 4'h1;
        10'd526: data = 4'h5;
        10'd527: data = 4'h6;
        10'd528: data = 4'h5;
        10'd529: data = 4'h0;
        10'd530: data = 4'h1;
        10'd531: data = 4'h1;
        10'd532: data = 4'h1;
        10'd533: data = 4'h5;
        10'd534: data = 4'h6;
        10'd535: data = 4'h6;
        10'd536: data = 4'h5;
        10'd537: data = 4'h5;
        10'd538: data = 4'h5;
        10'd539: data = 4'h5;
        10'd540: data = 4'h6;
        10'd541: data = 4'h6;
        10'd542: data = 4'h6;
        10'd543: data = 4'h5;
        10'd544: data = 4'h5;
        10'd545: data = 4'h5;
        10'd546: data = 4'h5;
        10'd547: data = 4'h6;
        10'd548: data = 4'h6;
        10'd549: data = 4'h6;
        10'd550: data = 4'h6;
        10'd551: data = 4'h6;
        10'd552: data = 4'h6;
        10'd553: data = 4'h6;
        10'd554: data = 4'h6;
        10'd555: data = 4'h6;
        10'd556: data = 4'h6;
        10'd557: data = 4'h6;
        10'd558: data = 4'h6;
        10'd559: data = 4'h6;
        10'd560: data = 4'h6;
        10'd561: data = 4'h6;
        10'd562: data = 4'h6;
        10'd563: data = 4'h6;
        10'd564: data = 4'h6;
        10'd565: data = 4'h6;
        10'd566: data = 4'h6;
        10'd567: data = 4'h6;
        10'd568: data = 4'h6;
        10'd569: data = 4'h6;
        10'd570: data = 4'h6;
        10'd571: data = 4'h6;
        10'd572: data = 4'h6;
        10'd573: data = 4'h6;
        10'd574: data = 4'h6;
        10'd575: data = 4'h6;
        10'd576: data = 4'h6;
        10'd577: data = 4'h6;
        10'd578: data = 4'h6;
        10'd579: data = 4'h6;
        10'd580: data = 4'h6;
        10'd581: data = 4'h6;
        10'd582: data = 4'h6;
        10'd583: data = 4'h6;
        10'd584: data = 4'h6;
        10'd585: data = 4'h6;
        10'd586: data = 4'h6;
        10'd587: data = 4'h6;
        10'd588: data = 4'h6;
        10'd589: data = 4'h6;
        10'd590: data = 4'h6;
        10'd591: data = 4'h6;
        10'd592: data = 4'h6;
        10'd593: data = 4'h6;
        10'd594: data = 4'h6;
        10'd595: data = 4'h6;
        10'd596: data = 4'h6;
        10'd597: data = 4'h6;
        10'd598: data = 4'h6;
        10'd599: data = 4'h6;
                10'd600: data = 4'h6;
        10'd601: data = 4'h6;
        10'd602: data = 4'h6;
        10'd603: data = 4'h6;
        10'd604: data = 4'h6;
        10'd605: data = 4'h6;
        10'd606: data = 4'h6;
        10'd607: data = 4'h6;
        10'd608: data = 4'h6;
        10'd609: data = 4'h6;
        10'd610: data = 4'h6;
        10'd611: data = 4'h6;
        10'd612: data = 4'h6;
        10'd613: data = 4'h6;
        10'd614: data = 4'h6;
        10'd615: data = 4'h6;
        10'd616: data = 4'h6;
        10'd617: data = 4'h6;
        10'd618: data = 4'h6;
        10'd619: data = 4'h6;
        10'd620: data = 4'h6;
        10'd621: data = 4'h6;
        10'd622: data = 4'h6;
        10'd623: data = 4'h6;
        10'd624: data = 4'h6;
        10'd625: data = 4'h6;
        10'd626: data = 4'h6;
        10'd627: data = 4'h6;
        10'd628: data = 4'h6;
        10'd629: data = 4'h6;
        10'd630: data = 4'h6;
        10'd631: data = 4'h6;
        10'd632: data = 4'h6;
        10'd633: data = 4'h6;
        10'd634: data = 4'h6;
        10'd635: data = 4'h6;
        10'd636: data = 4'h6;
        10'd637: data = 4'h6;
        10'd638: data = 4'h6;
        10'd639: data = 4'h6;
        default: data = 4'h0;
    endcase
end

endmodule


